`timescale 1 us / 100 ns
module har_front_end_tb();
	parameter inWidth = 15;
	parameter weightWidth = 16;
	parameter featureWidth = 16;
	//inputs
	logic clk;
	logic reset;
	logic weight_valid_NN;
	logic feature_valid_NN;
	logic signed [((inWidth-1)*weightWidth)-1:0] feature;
	logic signed [weightWidth-1:0] weight;
	//outputs
	logic output_valid_NN;
	logic [15:0] max_out_NN;
	logic [2:0] maxindex_out_NN;
	logic waiting_weight_NN;
	logic NN_busy;
	// wire signed [4*featureWidth-1:0] layer1Out;
	// wire signed [8*featureWidth-1:0] layer2Out;
	// wire signed [7*featureWidth-1:0] layer3Out;
	
	//read these from file
	
	logic signed [weightWidth-1:0] weightsL1[15*16-1:0]; // 224 weights for layer 1
	logic signed [weightWidth-1:0] weightsL2[17*16-1:0]; // 256 weights for layer 2
	logic signed [weightWidth-1:0] weightsL3[17*16-1:0]; // 256 weights for layer 3
	logic signed [weightWidth-1:0] weightsL4[17*3-1:0]; // 48 weights for layer 4
	integer f,i;
		
	initial $readmemh("finalweights1_new", weightsL1); // read from weights file
	initial $readmemh("finalweights2", weightsL2); // read from weights file
	initial $readmemh("finalweights3", weightsL3); // read from weights file
	initial $readmemh("finalweights4", weightsL4); // read from weights file
	//initial $readmemh("features", features); // read from features file
	
	har_front_end_logic_main  har_UUT (clk, reset, weight_valid_NN, feature_valid_NN, feature, weight, output_valid_NN, max_out_NN, maxindex_out_NN, NN_busy, waiting_weight_NN);
		
	//
	initial clk=0; //set up clock
	always #5 clk=~clk;
	
	/* initial begin
		//$fdumpfile("HAR_weight_load_wclockgate_100k.vcd");
		$fdumpvars (0, har_front_end_tb, "HAR_weight_load_wclockgate_100k.vcd");
		$fdumpon("HAR_weight_load_wclockgate_100k.vcd");
		#(6015) $fdumpoff("HAR_weight_load_wclockgate_100k.vcd");
		$fdumpflush("HAR_weight_load_wclockgate_100k.vcd");
	end
	
	initial begin
		#(6015) 
		//$fdumpfile("HAR_forward_mode_wclockgate_100k.vcd");
		$fdumpvars (0, har_front_end_tb,"HAR_forward_mode_wclockgate_100k.vcd");
		$fdumpon("HAR_forward_mode_wclockgate_100k.vcd");
		#(30000) $fdumpoff("HAR_forward_mode_wclockgate_100k.vcd");
		$fdumpflush("HAR_forward_mode_wclockgate_100k.vcd");
		$finish;
	end */

	initial begin
    f = $fopen("output.txt","w");

    for (i = 0; i<10000; i=i+1) begin
      @(posedge output_valid_NN);
      //$display("LFSR %b", out);
      $fwrite(f,"MAX:%d IDX:%d\n",   max_out_NN, maxindex_out_NN);
    end

    $fclose(f);  
    $finish;
  end
	
	initial begin // reset once
	reset=0;
	weight=0; 
	weight_valid_NN = 0;
	feature = 0;
	feature_valid_NN = 0;
	@(posedge clk)
	#1 reset=1;
	@(posedge clk)
	#1 reset=1;
	@(posedge clk)
	#1 reset=0;
	//weight loading
	@(posedge waiting_weight_NN)
			#1 weight_valid_NN = 1'b1;
			for(i=0;i<240;i=i+1) begin // write weights into the register
				@(posedge clk)
				#1 weight_valid_NN = 1'b1;
				#1 weight = weightsL1[i][15:0];
			end
			for(i=0;i<272;i=i+1) begin // write weights into the register
				@(posedge clk)
				#1 weight_valid_NN = 1'b1;
				#1 weight = weightsL2[i][15:0];
			end
	
			for(i=0;i<272;i=i+1) begin // write weights into the register
				@(posedge clk)
				#1 weight_valid_NN = 1'b1;
				#1 weight = weightsL3[i][15:0];
			end
			
			for(i=0;i<51;i=i+1) begin // write weights into the register
				@(posedge clk)
				#1 weight_valid_NN = 1'b1;
				#1 weight = weightsL4[i][15:0];
			end
		@(posedge clk);
	#1 weight_valid_NN = 1'b0;

	for(i=0;i<100;i=i+1) 
		@(posedge clk);
	//#10 feature = 224'b00000000000000000000000000000000000000000000000000000000000000100000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100; 
	#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010101000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010100110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010010010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001111011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001110111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000011010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000011010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000011000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000001000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000010100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000110011010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000110001010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000101101100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000101100100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000101111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001111000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001110000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001100001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001011101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100001000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000110100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000110010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000011110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000010110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000110111100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000001011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000010110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000010110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000001110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000011011010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000110000000011011001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000010000000011010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000001001100000000000000000000000011010110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000110011100000000011000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000110001100000000010111011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000101101110000000010101100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000101100110000000010101000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000011100100000000000010110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000010111000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010111011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010111001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010100101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010011101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000010101110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000100100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000011100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000011010011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000011001011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010111100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010111000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000001010010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001110101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001110011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001011111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001001000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100111010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000011100100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000011100000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000010111000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000010101000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000010001010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000010000010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000010100000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001110010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001110000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001011100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001010100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000110011100000000000101110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000110011000000000000101100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000101110000000000000011000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000101100000000000000010000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000101000010000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000001100000000101000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000100111010000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000100010000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000011011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000011010011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000011000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000011000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000001000010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000100000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000011110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000011010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000011110000000011000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000011010000000011000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000011100000000000000000000000010110011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000010000000010101100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000011100000000000000000000000010101011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000010000000000010100100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000011100000000000000000000000010011100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000001100000000000000000000000010011000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000110111100000000010010101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000110110100000000010010001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000101000000000000010010010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000011100000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000001000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000011000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000001010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000011100000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000011010001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000011001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000101000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000011011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000011010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010111010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010111000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010100100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010011100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000010110000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000110001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000101111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000010011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000110010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000110000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000011100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000010100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000111000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000100101000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000100100100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000011111100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000011101100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000011001110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000011000110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000001111110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000011010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000011000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000001000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000010100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000110011010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000110001010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000101101100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000101100100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000101111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001011010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001011000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000111100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000101101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000101001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000101110000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001101111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001101101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001011001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001010001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000111110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000101000110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001010100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001010010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000111110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000110110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000100111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000100011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000101111100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010110011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010110001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010011101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010010101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010000110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000010111110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000011110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000001000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000011011101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000011001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000011001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000101110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001101101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001100101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001010110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001010010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100011110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000110001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000101111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000010011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000011010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000011010000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000010101000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000010011000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000001111010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000001110010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000010101000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011011001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000011000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010111101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010101110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010101010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000001101110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001101000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001100110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001010010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000111011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000110111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000101010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001011000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001010110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000111010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000101011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000100111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000101110100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010110001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010101001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010011010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010010110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000010010110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000101000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000100010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000111010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000111000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000100100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000011100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000110110000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001011001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000111011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000101100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000101000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000101110010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000101101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000101011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000001111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010011101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001111111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001110000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001101100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000011101010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000010100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000010010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000010010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000010000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000001000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010011010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010011000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001111100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001101101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001101001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000100101110000000000011111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000100101010000000000011101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000100000010000000000001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000011110010000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000111000000000011110000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000011010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000011001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000001111011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010001011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001110111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001101111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001100000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001011100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100001010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000010000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000011011111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000011011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000100110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000100100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000010000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000001000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000001110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010010100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010010010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001111110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001110110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001100111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001100011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000011111100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010110110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010101110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010011111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000010001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011010110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011010100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000011000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010111000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010101001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010100101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000011101010000000000111001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000011100110000000000110111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000010111110000000000100011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000010101110000000000011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000010010000000000000001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000010001000000000000001000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000001101100100000000001111000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000001001110100000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011001011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010110111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010101111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010100000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010011100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000010001010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011001011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010110101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010101101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010011110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010011010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000010001110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000101010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000101000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000010100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001111110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001111100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001101000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001100000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001010001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100101000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001100101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001100010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001000110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000110111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000110011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000101011100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001111101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001111011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001100111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001011111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001010000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000101110100000000000100101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000101110000000000000100011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000101001000000000000001111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000001100000000100111110000000000001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000001000000000100111000000000000000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000101000000000100101010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000001000000000100011010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000100010110000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000001001000000000100010010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000011101110000000011001111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000011011110000000011000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000011000000000000010111000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000010111000000000010110100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000001000010100000000000000000000000001011000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000010110100000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000011011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000011010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000100101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000100011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000001111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000010000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010110100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010110001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010011101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010010101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010000110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000010111110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001111000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001110101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001100001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001011001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001000110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100110110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000111111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000101011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000100011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000010100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000010000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000110100010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000110011110000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000110011010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000101110010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000101100010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000101000100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000100111100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000001000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001101111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001101101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001011001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001010001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000111110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000101000110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001110001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001101001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001011010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001010110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100010110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010001011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001110111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001101111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001100000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001011100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100001010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001101010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001101000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001010100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000111101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000111001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000101010000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010101000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010100110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010010010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001111011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001110111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000011010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010101110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010101100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010011000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010010000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001111101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000101011010000000001001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000101010100000000001000110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000100101100000000000110010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000100011100000000000101010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000011111110000000000011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000011110110000000000010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000001100101000000000011001000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000110011000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001011110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001011100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000001100000000001001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000001000000000001001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000001000000000000000000000000000001001000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000100000000000000000000000000001000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000001110000000000111000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000100000000000000000000000000110001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000110000000000110000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000110000000000000000000000000000101101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000110101010000000000100001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000110100010000000000011101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000001100010000000000101101000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000001000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001100001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001011111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001001011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000110100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000110000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000101100010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000001011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000010110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000010110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000001110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000011011010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000011010110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000010110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000010001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010110110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010101110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010011111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000010001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011010101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000011000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010111001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010101010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010100110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000011111010000000001000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000011110100000000000111111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000011001100000000000101011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000010111100000000000100011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000010011110000000000010100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000010010110000000000010000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000001101000100000000001110110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000001001100000000000000000100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000001001011000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000001001011000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000001000001000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000111101000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000110101100000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000110011100000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000001111010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001111111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001111101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001101001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001100001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001010010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100100110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001101011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001101001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001010101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000111110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000111010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000110100010000000000101010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000110011110000000000101000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000101110110000000000010100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000101100110000000000001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000001100000000101001110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000101001000000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000101000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000001010100000000001101011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000001001110000000001101000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000100110000000001010100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000010110000000001001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000010000000000000000000000000001000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000111101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000111001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000101010000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001101011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001101001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001010101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000111110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000111010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000101001110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001110110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001110100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001100000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001011000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100111000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001110101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001110011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001011111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001001000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100111010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010101101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010101011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010001111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001111100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000011001010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010100100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010100010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010000110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001110111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001110011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000100110110000000000101101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000100110000000000000101010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000100001000000000000010110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000011111000000000000001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000100000000011011100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000011011010000000000000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000011010010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000001111000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000011111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000011101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000011100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010101010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010100111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010010011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010001011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001111100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001111000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000011010010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011100000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000011001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000011000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010110101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010110001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000001100000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000111101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000111011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000100111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000011111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000010000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000110101010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000100100010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000100011110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000011110110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000011100110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000011001000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000011000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000010000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001111011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001111001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001100101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001011101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100101110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000011111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000011101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000011100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001100101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001100011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001001111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000111000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000110100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000111000000000000000110011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000110111100000000000110001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000110010100000000000011101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000110000100000000000010101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000101100110000000000000110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000101011110000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000001101111100000000101011010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000001011011100000000100001010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000001011010000000000100000100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000001010000000000000011011100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000001001100000000000011001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000001000100100000000010101110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000001000010100000000010100110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000011001000000000000000000000000010001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000001011100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010110011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010110001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010011101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010010101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010000110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000010111110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000111010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000111000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000100100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000011100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000110110000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001110000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001101101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001011001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001010001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000111110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000101001100000000000000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000101001000000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000001001100000000101000110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000100100000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000100010000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000011110010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000011101010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000010010000000000010110100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000010001100000000010110010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000001100100000000010011110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000001010100000000010010110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000110110000000010000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000101110000000010000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000001100101000000000000000000000000001101100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000101111000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000011011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000011010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000100000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000011010001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000011001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010111010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010110110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000001010110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001010100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001010010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000111110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000110110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000100111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000100011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000101111100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000010010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000001110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000011011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000011010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001110000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001101110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001011010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001010010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000111111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000101000100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001101010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001101000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001010100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000111101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000111001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000101010000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011010000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010111010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010110010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010100011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010011111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000010000100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000110110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000101110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000011111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000110001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001111101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001101001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001100001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001010010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100100110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000011110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000010110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000011010110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000011001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010111111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010111011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000001001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000110000000000001000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000010000000000000110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000001001100000000000000000000000000000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000111000000000000010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000101000000000000001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000010000000000000000000000000011011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000011010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000010000000000011010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000001101100100000000000000000000000011001111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000001100101000000000000000000000000011000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000001100011000000000000000000000000010111100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000101000000000001001010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000110110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000101011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000101001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000010101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011001111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010111001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010110001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010100010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010011110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000110110110000000010011000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000110110010000000010010110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000110001010000000010000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000101111010000000001111010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000101011100000000001101011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000101010100000000001100111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000111101000000000010000110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000101001100000000000111000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000101000100000000000110100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000011110100000000000001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000011011100000000000000000000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000011010100000000000000100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000010011000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000010001000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000010111111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000011110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000001000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000011011101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000011001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000011001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000010100000000000000111001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000010011100000000000110111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000001110100000000000100011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000001100100000000000011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000001000110000000000001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000111110000000000001000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000001101111000000000000111000000000000000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000001101100100000000000101110000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000001101001100000000000100010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000001100001000000000000000000000000000000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000001011111100000000000000010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000001011011100000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000001010100000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000001010010000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000111101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011010001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011001111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010111011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010110011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010100100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010100000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000110001100000000010000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000110001000000000010000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000101100000000000001101111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000101010000000000001100111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000100110010000000001011000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000100101010000000001010100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000001000110100000000010000010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000100110000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000101100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000100100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000010101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000010001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000110100000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000011011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000011010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001100011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001100001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000110000000001001000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000010000000001000110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000001001100000000000000000000000001000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000010000000000000000000000000000110110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000110010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000010000000000000110010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000001101100100000000000000000000000000101010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000001100101000000000000000000000000000011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000001100011000000000000000000000000000010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000001010111100000000110010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000110110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000101110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000101100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000011000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000010000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010011101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010011010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010000110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001111110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000100000000001111110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000110100000000000000000000000001111100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000001110000000001101111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000110000000001101011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000001101111000000000000000000000000001101000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000001101011000000000000000000000000001100000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000001100011100000000000000000000000001010001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000001100001100000000000000000000000001001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000111011000000000100101000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000111100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010011101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001111111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001110000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001101100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000011101010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000010110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000001110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000011011010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000011010010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000011000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010111111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000001000100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010011001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010010110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001111010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001101011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001100111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000011110100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000011100100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000011100000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000010111000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000010101000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000010001010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000010000010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000010100000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001110101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001110011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001011111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001001000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100111010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010100110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010100100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010010000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010001000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001111001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001110101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000011011000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000010010010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000010001110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000001100110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000001010110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000111000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000110000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000011001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000100110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000010110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000001000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000001111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000110111010000000000001011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000110110110000000000001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000101100000000110100100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000011100000000110011100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000110001110000000011011010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000101111110000000011010010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000101100000000000011000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000101011000000000010111111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000011010100000000000000000000000000010011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000010001000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000011011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000011010011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000011000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000011000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000001000010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010110001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010101001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010011010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010010110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000010010110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011100000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000011001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000011000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010110101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010110001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000001100000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000101010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000100110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001010101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000111001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000101010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000100110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000101110110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000011010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010101100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010100100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010010101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010010001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000010100000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000110110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000101110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000011111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000110001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011011000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011010110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000011000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010111010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010101011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010100111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000100010100000000001010000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000100001110000000001001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000011100110000000000111001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000011010110000000000110001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000010111000000000000100010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000010110000000000000011110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000001100001100000000001110100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000001000100100000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000100111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000100101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000010001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001111111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001101011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001100011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001010100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001010000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100100010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001010001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001001111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000111011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000110011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000100100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000100000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000110000010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010110110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010101110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010011111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000010001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000111010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000111000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000100100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000011100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000110110000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001101111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001101101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001011001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000001000000000001010101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000010000000001010010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000001001100000000000000000000000001010001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000010000000000000000000000000001000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000111110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000010000000000000111110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000001101100100000000000000000000000000110110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000001100101000000000000000000000000000100111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000001100011000000000000000000000000000100011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000001010001100000000101111100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000110110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010100110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010100100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010010000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010001000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001111001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001110101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000011011000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001110110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001110100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001100000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001011000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100111000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000010010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000010000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000001000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000001000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000001011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000001000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000110111010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011011111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011011100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000011001000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000011000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010110001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010101101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000001101000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001011101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000111111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000110000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000101100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000101101010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010101100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010101010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010010110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001111111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001111011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000011001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000001011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000010010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000010010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000001010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000011011100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000011011000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000010010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010110110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010101110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010011111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000100000000000000000111010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000011111100000000000111000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000011010100000000000100100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000011000100000000000011100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000010100110000000000001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000010011110000000000001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000001101100000000000010001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000001001001000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000100110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010101011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010101000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010010100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001111101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001111001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000011010000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010000110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001110000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001101000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001011001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001010101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100011000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000011010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000110111100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000110101100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000110001110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000110000110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000011110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000011001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000010110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000101101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000101011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000001111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000101110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000100110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000010011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000110011100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000001110010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000001101110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000001000110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000110110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000011000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000010000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000011011001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000100100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000011100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000011010011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000011001111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000100100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000101001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000100111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000010011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000001011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000001000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000100000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000010000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000011000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000011010101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000011010001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000100000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001101110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001100110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001010011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100011100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010110011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010101011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010011100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010011000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000010010010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011001000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010110100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010101100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010011101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010011001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000010010000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010011101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001111111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001110000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001101100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000011101010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001110101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001110011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001011111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001001000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100111010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011010011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011010001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010111101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010110101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010100110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010100010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000001111110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010011000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010010101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001111001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001101010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001100110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000011110110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010000110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001110010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001101010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100010100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000100100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000011100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000011010011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000011001011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010111100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010111000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000001010010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010111010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010111000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010100100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010011100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010001101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010001001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000010110000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000101110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000101100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000011000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000010000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000001101000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000001100100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000111100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000101100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000001110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000011011110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000010010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000110011110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000110001110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000101110000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000101101000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000100101010000000011000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000100100110000000011000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000011111110000000010101100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000011101110000000010100100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000011010000000000010010101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000011001000000000010010001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000111110100000000000000000000000000101101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000101000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000010010111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000010010101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001111001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001101010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001100110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000011110110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011001010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010110110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010101110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010011111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000010001100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000100010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000011010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000110111100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000110101100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000110001110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000110000110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000011110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000011100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000001110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000011011110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000011001111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000011001011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000101100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000111000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000110000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000100001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000011101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000110001000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001111111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000001111101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000001101001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000001100001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000001010010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000001001110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000100100110000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000011000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000011000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000010101100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000010100100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000010010101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000010010001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000110100100000000010000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000110100000000000010000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000001000000000101111100000000001101110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000001000000000101111000000000001101100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000001000000000101101000000000001100100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000001000000000101001010000000001010101;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000001000000000101000010000000001010001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000001001001000000000010100000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000100001000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000001000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000010000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000110100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000110010;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000011110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000010110;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000110111100000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000111001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000110111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000100011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000011011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000001100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000001000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000110110010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000001000001;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000111111;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000101011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000100011;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000010100;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000010000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000110100010000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000001000000000110010000000000011001000000000001100100000000000110010000000000000001010000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000001100100000000000110010000000000011001000000000000000010000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000000000000000010100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000010000000000001000000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000100000000000001111000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000000110000000000000100000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;
#990 feature = 224'b00000000011001000000000001100100000000000110010000000000011001000000000000000000000000000110010000000000011001000000000001100100000000000110010000000000000001000000000011100001000000000000000000000000000000000000000000000000;
feature_valid_NN = 1'b1;
#10 feature_valid_NN = 1'b0;

	for(i=0;i<500;i=i+1) 
		@(posedge clk);
	
	//$fclose(filehandle);
	$finish;
end

endmodule